VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO logicfunctions
  CLASS BLOCK ;
  FOREIGN logicfunctions ;
  ORIGIN 2.600 0.000 ;
  SIZE 33.100 BY 13.100 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 1.400 0.800 1.800 4.500 ;
        RECT 3.800 0.800 4.200 4.500 ;
        RECT 6.200 0.800 6.600 3.100 ;
        RECT 8.600 0.800 9.000 3.100 ;
        RECT 10.200 0.800 10.600 3.100 ;
        RECT 11.800 0.800 12.200 4.500 ;
        RECT 14.200 0.800 14.600 3.100 ;
        RECT 15.000 0.800 15.400 3.100 ;
        RECT 16.600 0.800 17.000 5.100 ;
        RECT 19.800 0.800 20.200 5.100 ;
        RECT 23.000 0.800 23.400 4.500 ;
        RECT 27.000 0.800 27.400 3.100 ;
        RECT 0.200 0.200 27.800 0.800 ;
      LAYER via1 ;
        RECT 6.600 0.300 7.000 0.700 ;
        RECT 7.300 0.300 7.700 0.700 ;
      LAYER metal2 ;
        RECT 6.400 0.300 8.000 0.700 ;
      LAYER via2 ;
        RECT 6.600 0.300 7.000 0.700 ;
        RECT 7.300 0.300 7.700 0.700 ;
      LAYER metal3 ;
        RECT 6.400 0.300 8.000 0.700 ;
      LAYER via3 ;
        RECT 6.600 0.300 7.000 0.700 ;
        RECT 7.400 0.300 7.800 0.700 ;
      LAYER metal4 ;
        RECT 6.400 0.300 8.000 0.700 ;
      LAYER via4 ;
        RECT 6.600 0.300 7.000 0.700 ;
        RECT 7.300 0.300 7.700 0.700 ;
      LAYER metal5 ;
        RECT 6.400 0.200 8.000 0.700 ;
      LAYER via5 ;
        RECT 7.400 0.200 7.900 0.700 ;
      LAYER metal6 ;
        RECT 6.400 0.000 8.000 13.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.200 10.200 27.800 10.800 ;
        RECT 1.400 7.900 1.800 10.200 ;
        RECT 3.800 7.900 4.200 10.200 ;
        RECT 6.200 8.900 6.600 10.200 ;
        RECT 8.600 7.900 9.000 10.200 ;
        RECT 11.800 7.900 12.200 10.200 ;
        RECT 14.200 8.900 14.600 10.200 ;
        RECT 15.000 8.900 15.400 10.200 ;
        RECT 17.400 8.300 17.800 10.200 ;
        RECT 22.400 7.900 22.800 10.200 ;
        RECT 25.400 7.900 25.800 10.200 ;
        RECT 27.000 8.900 27.400 10.200 ;
      LAYER via1 ;
        RECT 20.200 10.300 20.600 10.700 ;
        RECT 20.900 10.300 21.300 10.700 ;
      LAYER metal2 ;
        RECT 20.000 10.300 21.600 10.700 ;
      LAYER via2 ;
        RECT 20.200 10.300 20.600 10.700 ;
        RECT 20.900 10.300 21.300 10.700 ;
      LAYER metal3 ;
        RECT 20.000 10.300 21.600 10.700 ;
      LAYER via3 ;
        RECT 20.200 10.300 20.600 10.700 ;
        RECT 21.000 10.300 21.400 10.700 ;
      LAYER metal4 ;
        RECT 20.000 10.300 21.600 10.700 ;
      LAYER via4 ;
        RECT 20.200 10.300 20.600 10.700 ;
        RECT 20.900 10.300 21.300 10.700 ;
      LAYER metal5 ;
        RECT 20.000 10.200 21.600 10.700 ;
      LAYER via5 ;
        RECT 21.000 10.200 21.500 10.700 ;
      LAYER metal6 ;
        RECT 20.000 0.000 21.600 13.000 ;
    END
  END gnd
  PIN x1
    PORT
      LAYER metal1 ;
        RECT 17.400 5.800 17.800 6.600 ;
        RECT 22.200 6.100 22.600 6.200 ;
        RECT 22.200 5.800 23.000 6.100 ;
        RECT 22.600 5.600 23.000 5.800 ;
      LAYER metal2 ;
        RECT 17.400 6.200 17.700 13.100 ;
        RECT 17.400 5.800 17.800 6.200 ;
        RECT 21.400 6.100 21.800 6.200 ;
        RECT 22.200 6.100 22.600 6.200 ;
        RECT 21.400 5.800 22.600 6.100 ;
      LAYER metal3 ;
        RECT 17.400 6.100 17.800 6.200 ;
        RECT 21.400 6.100 21.800 6.200 ;
        RECT 17.400 5.800 21.800 6.100 ;
    END
  END x1
  PIN x2
    PORT
      LAYER metal1 ;
        RECT 27.000 7.800 27.400 8.600 ;
        RECT 27.000 7.200 27.300 7.800 ;
        RECT 24.600 6.800 25.000 7.200 ;
        RECT 27.000 6.800 27.400 7.200 ;
        RECT 24.600 6.600 24.900 6.800 ;
        RECT 24.500 6.200 24.900 6.600 ;
      LAYER metal2 ;
        RECT 24.600 7.800 25.000 8.200 ;
        RECT 27.000 7.800 27.400 8.200 ;
        RECT 24.600 7.200 24.900 7.800 ;
        RECT 27.000 7.200 27.300 7.800 ;
        RECT 24.600 6.800 25.000 7.200 ;
        RECT 27.000 6.800 27.400 7.200 ;
      LAYER metal3 ;
        RECT 24.600 8.100 25.000 8.200 ;
        RECT 27.000 8.100 27.400 8.200 ;
        RECT 24.600 7.800 30.500 8.100 ;
    END
  END x2
  PIN x3
    PORT
      LAYER metal1 ;
        RECT 15.000 7.800 15.400 8.600 ;
        RECT 20.600 7.100 21.000 7.200 ;
        RECT 23.000 7.100 23.400 7.200 ;
        RECT 20.600 6.800 23.400 7.100 ;
        RECT 23.000 6.400 23.400 6.800 ;
      LAYER metal2 ;
        RECT 15.000 9.200 15.300 13.100 ;
        RECT 15.000 8.800 15.400 9.200 ;
        RECT 20.600 8.800 21.000 9.200 ;
        RECT 15.000 8.200 15.300 8.800 ;
        RECT 15.000 7.800 15.400 8.200 ;
        RECT 20.600 7.200 20.900 8.800 ;
        RECT 20.600 6.800 21.000 7.200 ;
      LAYER metal3 ;
        RECT 15.000 9.100 15.400 9.200 ;
        RECT 20.600 9.100 21.000 9.200 ;
        RECT 15.000 8.800 21.000 9.100 ;
    END
  END x3
  PIN x4
    PORT
      LAYER metal1 ;
        RECT 19.800 6.100 20.200 7.200 ;
        RECT 20.600 6.100 21.000 6.200 ;
        RECT 19.800 5.800 21.000 6.100 ;
        RECT 25.400 5.400 25.800 6.200 ;
      LAYER via1 ;
        RECT 20.600 5.800 21.000 6.200 ;
        RECT 25.400 5.800 25.800 6.200 ;
      LAYER metal2 ;
        RECT 20.600 5.800 21.000 6.200 ;
        RECT 25.400 5.800 25.800 6.200 ;
        RECT 20.600 5.200 20.900 5.800 ;
        RECT 25.400 5.200 25.700 5.800 ;
        RECT 20.600 4.800 21.000 5.200 ;
        RECT 25.400 4.800 25.800 5.200 ;
      LAYER metal3 ;
        RECT 25.400 6.100 25.800 6.200 ;
        RECT 25.400 5.800 30.500 6.100 ;
        RECT 20.600 5.100 21.000 5.200 ;
        RECT 25.400 5.100 25.800 5.200 ;
        RECT 20.600 4.800 25.800 5.100 ;
    END
  END x4
  PIN g
    PORT
      LAYER metal1 ;
        RECT 0.600 6.200 1.000 9.900 ;
        RECT 0.600 5.100 0.900 6.200 ;
        RECT 0.600 1.100 1.000 5.100 ;
      LAYER via1 ;
        RECT 0.600 6.800 1.000 7.200 ;
      LAYER metal2 ;
        RECT 0.600 6.800 1.000 7.200 ;
        RECT 0.600 6.200 0.900 6.800 ;
        RECT 0.600 5.800 1.000 6.200 ;
      LAYER metal3 ;
        RECT 0.600 6.100 1.000 6.200 ;
        RECT -2.600 5.800 1.000 6.100 ;
    END
  END g
  PIN h
    PORT
      LAYER metal1 ;
        RECT 11.000 6.200 11.400 9.900 ;
        RECT 11.000 5.100 11.300 6.200 ;
        RECT 11.000 1.100 11.400 5.100 ;
      LAYER via1 ;
        RECT 11.000 8.800 11.400 9.200 ;
      LAYER metal2 ;
        RECT 9.400 10.200 9.700 13.100 ;
        RECT 9.400 9.800 9.800 10.200 ;
        RECT 11.000 9.800 11.400 10.200 ;
        RECT 11.000 9.200 11.300 9.800 ;
        RECT 11.000 8.800 11.400 9.200 ;
      LAYER metal3 ;
        RECT 9.400 10.100 9.800 10.200 ;
        RECT 11.000 10.100 11.400 10.200 ;
        RECT 9.400 9.800 11.400 10.100 ;
    END
  END h
  PIN f
    PORT
      LAYER metal1 ;
        RECT 3.000 6.200 3.400 9.900 ;
        RECT 3.000 5.100 3.300 6.200 ;
        RECT 3.000 1.100 3.400 5.100 ;
      LAYER via1 ;
        RECT 3.000 7.800 3.400 8.200 ;
      LAYER metal2 ;
        RECT 3.000 8.800 3.400 9.200 ;
        RECT 3.000 8.200 3.300 8.800 ;
        RECT 3.000 7.800 3.400 8.200 ;
      LAYER metal3 ;
        RECT 3.000 8.800 3.400 9.200 ;
        RECT 3.000 8.100 3.300 8.800 ;
        RECT -2.600 7.800 3.300 8.100 ;
    END
  END f
  OBS
      LAYER metal1 ;
        RECT 2.200 7.600 2.600 9.900 ;
        RECT 4.600 7.600 5.000 9.900 ;
        RECT 1.500 7.300 2.600 7.600 ;
        RECT 3.900 7.300 5.000 7.600 ;
        RECT 1.500 5.800 1.800 7.300 ;
        RECT 2.200 5.800 2.600 6.600 ;
        RECT 3.900 5.800 4.200 7.300 ;
        RECT 4.600 5.800 5.000 6.600 ;
        RECT 1.200 5.400 1.800 5.800 ;
        RECT 3.600 5.400 4.200 5.800 ;
        RECT 1.500 5.100 1.800 5.400 ;
        RECT 3.900 5.100 4.200 5.400 ;
        RECT 1.500 4.800 2.600 5.100 ;
        RECT 3.900 4.800 5.000 5.100 ;
        RECT 2.200 1.100 2.600 4.800 ;
        RECT 4.600 1.100 5.000 4.800 ;
        RECT 5.400 1.100 5.800 9.900 ;
        RECT 6.200 7.800 6.600 8.600 ;
        RECT 9.900 8.200 10.300 9.900 ;
        RECT 9.400 7.900 10.300 8.200 ;
        RECT 6.200 7.100 6.500 7.800 ;
        RECT 8.600 7.100 9.000 7.600 ;
        RECT 6.200 6.800 9.000 7.100 ;
        RECT 8.600 6.200 8.900 6.800 ;
        RECT 8.600 5.800 9.000 6.200 ;
        RECT 9.400 6.100 9.800 7.900 ;
        RECT 12.600 7.600 13.000 9.900 ;
        RECT 11.900 7.300 13.000 7.600 ;
        RECT 10.200 6.100 10.600 6.200 ;
        RECT 9.400 5.800 10.600 6.100 ;
        RECT 11.900 5.800 12.200 7.300 ;
        RECT 12.600 6.100 13.000 6.600 ;
        RECT 13.400 6.100 13.800 9.900 ;
        RECT 14.200 7.800 14.600 8.600 ;
        RECT 12.600 5.800 13.800 6.100 ;
        RECT 9.400 1.100 9.800 5.800 ;
        RECT 11.600 5.400 12.200 5.800 ;
        RECT 10.200 4.400 10.600 5.200 ;
        RECT 11.900 5.100 12.200 5.400 ;
        RECT 11.900 4.800 13.000 5.100 ;
        RECT 12.600 1.100 13.000 4.800 ;
        RECT 13.400 1.100 13.800 5.800 ;
        RECT 15.800 7.100 16.200 9.900 ;
        RECT 16.600 8.000 17.000 9.900 ;
        RECT 18.200 9.600 20.200 9.900 ;
        RECT 18.200 8.000 18.600 9.600 ;
        RECT 16.600 7.900 18.600 8.000 ;
        RECT 19.000 7.900 19.400 9.300 ;
        RECT 19.800 7.900 20.200 9.600 ;
        RECT 23.700 7.900 24.500 9.900 ;
        RECT 16.700 7.700 18.500 7.900 ;
        RECT 17.000 7.200 17.400 7.400 ;
        RECT 19.100 7.200 19.400 7.900 ;
        RECT 23.900 7.200 24.200 7.900 ;
        RECT 16.600 7.100 17.400 7.200 ;
        RECT 15.800 6.900 17.400 7.100 ;
        RECT 18.200 6.900 19.400 7.200 ;
        RECT 15.800 6.800 17.000 6.900 ;
        RECT 18.200 6.800 18.600 6.900 ;
        RECT 23.800 6.800 24.200 7.200 ;
        RECT 15.800 1.100 16.200 6.800 ;
        RECT 18.200 5.100 18.500 6.800 ;
        RECT 19.000 5.800 19.400 6.600 ;
        RECT 23.900 6.200 24.200 6.800 ;
        RECT 23.800 5.800 24.200 6.200 ;
        RECT 23.900 5.700 24.200 5.800 ;
        RECT 23.900 5.400 24.900 5.700 ;
        RECT 24.600 5.100 24.900 5.400 ;
        RECT 17.900 1.100 18.900 5.100 ;
        RECT 22.200 4.800 24.200 5.100 ;
        RECT 22.200 1.100 22.600 4.800 ;
        RECT 23.800 1.400 24.200 4.800 ;
        RECT 24.600 1.700 25.000 5.100 ;
        RECT 25.400 1.400 25.800 5.100 ;
        RECT 23.800 1.100 25.800 1.400 ;
        RECT 26.200 1.100 26.600 9.900 ;
      LAYER via1 ;
        RECT 5.400 6.800 5.800 7.200 ;
        RECT 10.200 5.800 10.600 6.200 ;
        RECT 10.200 4.800 10.600 5.200 ;
        RECT 26.200 8.800 26.600 9.200 ;
      LAYER metal2 ;
        RECT 26.200 9.100 26.600 9.200 ;
        RECT 27.000 9.100 27.400 9.200 ;
        RECT 26.200 8.800 27.400 9.100 ;
        RECT 13.400 8.100 13.800 8.200 ;
        RECT 14.200 8.100 14.600 8.200 ;
        RECT 13.400 7.800 14.600 8.100 ;
        RECT 18.200 7.800 18.600 8.200 ;
        RECT 19.000 7.800 19.400 8.200 ;
        RECT 2.200 6.800 2.600 7.200 ;
        RECT 4.600 7.100 5.000 7.200 ;
        RECT 5.400 7.100 5.800 7.200 ;
        RECT 4.600 6.800 5.800 7.100 ;
        RECT 8.600 6.800 9.000 7.200 ;
        RECT 2.200 6.200 2.500 6.800 ;
        RECT 8.600 6.200 8.900 6.800 ;
        RECT 2.200 5.800 2.600 6.200 ;
        RECT 4.600 6.100 5.000 6.200 ;
        RECT 5.400 6.100 5.800 6.200 ;
        RECT 4.600 5.800 5.800 6.100 ;
        RECT 8.600 5.800 9.000 6.200 ;
        RECT 9.400 6.100 9.800 6.200 ;
        RECT 10.200 6.100 10.600 6.200 ;
        RECT 9.400 5.800 10.600 6.100 ;
        RECT 13.400 5.200 13.700 7.800 ;
        RECT 18.200 7.200 18.500 7.800 ;
        RECT 18.200 6.800 18.600 7.200 ;
        RECT 19.000 6.200 19.300 7.800 ;
        RECT 23.000 7.100 23.400 7.200 ;
        RECT 23.800 7.100 24.200 7.200 ;
        RECT 23.000 6.800 24.200 7.100 ;
        RECT 19.000 5.800 19.400 6.200 ;
        RECT 10.200 5.100 10.600 5.200 ;
        RECT 11.000 5.100 11.400 5.200 ;
        RECT 10.200 4.800 11.400 5.100 ;
        RECT 13.400 4.800 13.800 5.200 ;
      LAYER via2 ;
        RECT 27.000 8.800 27.400 9.200 ;
        RECT 5.400 5.800 5.800 6.200 ;
        RECT 11.000 4.800 11.400 5.200 ;
      LAYER metal3 ;
        RECT 27.000 9.100 27.400 9.200 ;
        RECT 21.400 8.800 27.400 9.100 ;
        RECT 13.400 8.100 13.800 8.200 ;
        RECT 18.200 8.100 18.600 8.200 ;
        RECT 13.400 7.800 18.600 8.100 ;
        RECT 19.000 8.100 19.400 8.200 ;
        RECT 21.400 8.100 21.700 8.800 ;
        RECT 19.000 7.800 21.700 8.100 ;
        RECT 2.200 7.100 2.600 7.200 ;
        RECT 4.600 7.100 5.000 7.200 ;
        RECT 2.200 6.800 5.000 7.100 ;
        RECT 8.600 7.100 9.000 7.200 ;
        RECT 23.000 7.100 23.400 7.200 ;
        RECT 8.600 6.800 23.400 7.100 ;
        RECT 5.400 6.100 5.800 6.200 ;
        RECT 9.400 6.100 9.800 6.200 ;
        RECT 5.400 5.800 9.800 6.100 ;
        RECT 11.000 5.100 11.400 5.200 ;
        RECT 13.400 5.100 13.800 5.200 ;
        RECT 11.000 4.800 13.800 5.100 ;
  END
END logicfunctions
END LIBRARY

