* NGSPICE file created from boolean_equation.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

.subckt boolean_equation vdd gnd A B C D E F
XFILL_0_0_0 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XNAND3X1_1 D C E gnd AND2X2_1/A vdd NAND3X1
XBUFX2_1 BUFX2_1/A gnd F vdd BUFX2
XNAND2X1_1 B A gnd AND2X2_1/B vdd NAND2X1
XFILL_0_1_0 gnd vdd FILL
XFILL_0_1_1 gnd vdd FILL
XAND2X2_1 AND2X2_1/A AND2X2_1/B gnd BUFX2_1/A vdd AND2X2
.ends

