VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO boolean_equation
  CLASS BLOCK ;
  FOREIGN boolean_equation ;
  ORIGIN 2.600 0.000 ;
  SIZE 20.300 BY 11.000 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.800 1.000 3.100 ;
        RECT 2.200 0.800 2.600 3.100 ;
        RECT 5.400 0.800 5.800 4.500 ;
        RECT 7.800 0.800 8.200 4.900 ;
        RECT 9.400 0.800 9.800 3.100 ;
        RECT 12.600 0.800 13.000 2.900 ;
        RECT 14.200 0.800 14.600 3.100 ;
        RECT 0.200 0.200 15.000 0.800 ;
      LAYER via1 ;
        RECT 2.600 0.300 3.000 0.700 ;
        RECT 3.300 0.300 3.700 0.700 ;
      LAYER metal2 ;
        RECT 2.400 0.300 4.000 0.700 ;
      LAYER via2 ;
        RECT 2.600 0.300 3.000 0.700 ;
        RECT 3.300 0.300 3.700 0.700 ;
      LAYER metal3 ;
        RECT 2.400 0.300 4.000 0.700 ;
      LAYER via3 ;
        RECT 2.600 0.300 3.000 0.700 ;
        RECT 3.400 0.300 3.800 0.700 ;
      LAYER metal4 ;
        RECT 2.400 0.300 4.000 0.700 ;
      LAYER via4 ;
        RECT 2.600 0.300 3.000 0.700 ;
        RECT 3.300 0.300 3.700 0.700 ;
      LAYER metal5 ;
        RECT 2.400 0.200 4.000 0.700 ;
      LAYER via5 ;
        RECT 3.400 0.200 3.900 0.700 ;
      LAYER metal6 ;
        RECT 2.400 0.000 4.000 11.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.200 10.200 15.000 10.800 ;
        RECT 0.600 7.900 1.000 10.200 ;
        RECT 5.400 7.900 5.800 10.200 ;
        RECT 8.100 8.000 8.500 10.200 ;
        RECT 14.200 6.900 14.600 10.200 ;
      LAYER via1 ;
        RECT 9.800 10.300 10.200 10.700 ;
        RECT 10.500 10.300 10.900 10.700 ;
      LAYER metal2 ;
        RECT 9.600 10.300 11.200 10.700 ;
      LAYER via2 ;
        RECT 9.800 10.300 10.200 10.700 ;
        RECT 10.500 10.300 10.900 10.700 ;
      LAYER metal3 ;
        RECT 9.600 10.300 11.200 10.700 ;
      LAYER via3 ;
        RECT 9.800 10.300 10.200 10.700 ;
        RECT 10.600 10.300 11.000 10.700 ;
      LAYER metal4 ;
        RECT 9.600 10.300 11.200 10.700 ;
      LAYER via4 ;
        RECT 9.800 10.300 10.200 10.700 ;
        RECT 10.500 10.300 10.900 10.700 ;
      LAYER metal5 ;
        RECT 9.600 10.200 11.200 10.700 ;
      LAYER via5 ;
        RECT 10.600 10.200 11.100 10.700 ;
      LAYER metal6 ;
        RECT 9.600 0.000 11.200 11.000 ;
    END
  END gnd
  PIN A
    PORT
      LAYER metal1 ;
        RECT 2.200 4.400 2.600 5.200 ;
      LAYER via1 ;
        RECT 2.200 4.800 2.600 5.200 ;
      LAYER metal2 ;
        RECT 2.200 5.800 2.600 6.200 ;
        RECT 2.200 5.200 2.500 5.800 ;
        RECT 2.200 4.800 2.600 5.200 ;
      LAYER metal3 ;
        RECT 2.200 6.100 2.600 6.200 ;
        RECT -2.600 5.800 2.600 6.100 ;
    END
  END A
  PIN B
    PORT
      LAYER metal1 ;
        RECT 0.600 6.800 1.000 7.600 ;
      LAYER metal2 ;
        RECT 0.600 9.800 1.000 10.200 ;
        RECT 0.600 7.200 0.900 9.800 ;
        RECT 0.600 6.800 1.000 7.200 ;
      LAYER metal3 ;
        RECT 0.600 10.100 1.000 10.200 ;
        RECT -2.600 9.800 1.000 10.100 ;
    END
  END B
  PIN C
    PORT
      LAYER metal1 ;
        RECT 13.000 5.800 13.800 6.200 ;
      LAYER via1 ;
        RECT 13.400 5.800 13.800 6.200 ;
      LAYER metal2 ;
        RECT 13.400 7.800 13.800 8.200 ;
        RECT 13.400 6.200 13.700 7.800 ;
        RECT 13.400 5.800 13.800 6.200 ;
      LAYER metal3 ;
        RECT 13.400 8.100 13.800 8.200 ;
        RECT 13.400 7.800 17.700 8.100 ;
    END
  END C
  PIN D
    PORT
      LAYER metal1 ;
        RECT 14.200 4.800 14.600 6.200 ;
      LAYER via1 ;
        RECT 14.200 5.800 14.600 6.200 ;
      LAYER metal2 ;
        RECT 14.200 5.800 14.600 6.200 ;
        RECT 14.200 5.200 14.500 5.800 ;
        RECT 14.200 4.800 14.600 5.200 ;
      LAYER metal3 ;
        RECT 14.200 5.800 17.700 6.100 ;
        RECT 14.200 5.200 14.500 5.800 ;
        RECT 14.200 4.800 14.600 5.200 ;
    END
  END D
  PIN E
    PORT
      LAYER metal1 ;
        RECT 12.600 4.100 13.000 4.600 ;
        RECT 13.400 4.100 13.800 4.200 ;
        RECT 12.600 3.800 13.800 4.100 ;
      LAYER via1 ;
        RECT 13.400 3.800 13.800 4.200 ;
      LAYER metal2 ;
        RECT 13.400 4.100 13.800 4.200 ;
        RECT 14.200 4.100 14.600 4.200 ;
        RECT 13.400 3.800 14.600 4.100 ;
      LAYER via2 ;
        RECT 14.200 3.800 14.600 4.200 ;
      LAYER metal3 ;
        RECT 14.200 4.100 14.600 4.200 ;
        RECT 14.200 3.800 17.700 4.100 ;
    END
  END E
  PIN F
    PORT
      LAYER metal1 ;
        RECT 3.800 8.100 4.200 8.200 ;
        RECT 4.600 8.100 5.000 9.900 ;
        RECT 3.800 7.800 5.000 8.100 ;
        RECT 4.600 6.200 5.000 7.800 ;
        RECT 4.600 5.100 4.900 6.200 ;
        RECT 4.600 1.100 5.000 5.100 ;
      LAYER metal2 ;
        RECT 3.000 8.100 3.400 8.200 ;
        RECT 3.800 8.100 4.200 8.200 ;
        RECT 3.000 7.800 4.200 8.100 ;
      LAYER metal3 ;
        RECT 3.000 8.100 3.400 8.200 ;
        RECT -2.600 7.800 3.400 8.100 ;
    END
  END F
  OBS
      LAYER metal1 ;
        RECT 1.900 8.200 2.300 9.900 ;
        RECT 1.400 7.900 2.300 8.200 ;
        RECT 1.400 7.100 1.800 7.900 ;
        RECT 6.200 7.600 6.600 9.900 ;
        RECT 7.300 8.400 7.700 9.900 ;
        RECT 5.500 7.300 6.600 7.600 ;
        RECT 7.000 7.900 7.700 8.400 ;
        RECT 9.400 7.900 9.800 9.900 ;
        RECT 3.000 7.100 3.400 7.200 ;
        RECT 1.400 6.800 3.400 7.100 ;
        RECT 1.400 1.100 1.800 6.800 ;
        RECT 5.500 5.800 5.800 7.300 ;
        RECT 6.200 6.100 6.600 6.600 ;
        RECT 7.000 6.200 7.300 7.900 ;
        RECT 9.400 7.800 9.700 7.900 ;
        RECT 8.800 7.600 9.700 7.800 ;
        RECT 7.600 7.500 9.700 7.600 ;
        RECT 7.600 7.300 9.100 7.500 ;
        RECT 7.600 7.200 8.000 7.300 ;
        RECT 7.000 6.100 7.400 6.200 ;
        RECT 6.200 5.800 7.400 6.100 ;
        RECT 5.200 5.400 5.800 5.800 ;
        RECT 5.500 5.100 5.800 5.400 ;
        RECT 7.000 5.100 7.300 5.800 ;
        RECT 7.700 5.500 8.000 7.200 ;
        RECT 9.400 7.100 9.800 7.200 ;
        RECT 12.400 7.100 12.800 9.900 ;
        RECT 8.400 6.600 9.000 7.000 ;
        RECT 9.400 6.900 12.800 7.100 ;
        RECT 9.400 6.800 12.700 6.900 ;
        RECT 8.600 6.200 8.900 6.600 ;
        RECT 9.400 6.400 9.800 6.800 ;
        RECT 8.600 5.800 9.000 6.200 ;
        RECT 7.700 5.200 8.900 5.500 ;
        RECT 11.900 5.200 12.200 6.800 ;
        RECT 5.500 4.800 6.600 5.100 ;
        RECT 6.200 1.100 6.600 4.800 ;
        RECT 7.000 1.100 7.400 5.100 ;
        RECT 8.600 3.100 8.900 5.200 ;
        RECT 11.800 4.800 12.200 5.200 ;
        RECT 11.900 3.500 12.200 4.800 ;
        RECT 11.900 3.200 13.700 3.500 ;
        RECT 11.900 3.100 12.200 3.200 ;
        RECT 8.600 1.100 9.000 3.100 ;
        RECT 11.800 1.100 12.200 3.100 ;
        RECT 13.400 3.100 13.700 3.200 ;
        RECT 13.400 1.100 13.800 3.100 ;
      LAYER via1 ;
        RECT 3.000 6.800 3.400 7.200 ;
        RECT 8.600 6.600 9.000 7.000 ;
      LAYER metal2 ;
        RECT 3.000 7.100 3.400 7.200 ;
        RECT 3.800 7.100 4.200 7.200 ;
        RECT 3.000 6.800 4.200 7.100 ;
        RECT 7.800 6.900 8.200 7.000 ;
        RECT 8.600 6.900 9.000 7.000 ;
        RECT 7.800 6.600 9.000 6.900 ;
      LAYER via2 ;
        RECT 3.800 6.800 4.200 7.200 ;
      LAYER metal3 ;
        RECT 3.800 7.100 4.200 7.200 ;
        RECT 3.800 7.000 8.100 7.100 ;
        RECT 3.800 6.800 8.200 7.000 ;
        RECT 7.800 6.600 8.200 6.800 ;
  END
END boolean_equation
END LIBRARY

