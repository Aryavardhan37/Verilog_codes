* NGSPICE file created from logicfunctions.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

.subckt logicfunctions vdd gnd x1 x2 x3 x4 g h f
XFILL_0_0_0 gnd vdd FILL
XAOI22X1_1 x1 x3 x4 x2 gnd INVX1_3/A vdd AOI22X1
XFILL_0_0_1 gnd vdd FILL
XBUFX2_1 BUFX2_1/A gnd f vdd BUFX2
XBUFX2_2 BUFX2_2/A gnd g vdd BUFX2
XBUFX2_3 BUFX2_3/A gnd h vdd BUFX2
XFILL_0_1_0 gnd vdd FILL
XNAND2X1_1 INVX1_3/A INVX1_2/A gnd BUFX2_1/A vdd NAND2X1
XFILL_0_1_1 gnd vdd FILL
XINVX1_1 x2 gnd INVX1_1/Y vdd INVX1
XINVX1_2 INVX1_2/A gnd BUFX2_3/A vdd INVX1
XOAI22X1_1 INVX1_4/Y x1 x4 INVX1_1/Y gnd INVX1_2/A vdd OAI22X1
XINVX1_3 INVX1_3/A gnd BUFX2_2/A vdd INVX1
XINVX1_4 x3 gnd INVX1_4/Y vdd INVX1
.ends

