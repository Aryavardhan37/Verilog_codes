VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO full_adder
  CLASS BLOCK ;
  FOREIGN full_adder ;
  ORIGIN 1.900 0.000 ;
  SIZE 19.900 BY 24.000 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 7.600 1.600 8.400 9.000 ;
        RECT 12.400 1.600 13.200 9.000 ;
        RECT 0.400 0.400 15.600 1.600 ;
      LAYER via1 ;
        RECT 1.600 0.800 2.000 1.200 ;
        RECT 3.000 0.800 3.400 1.200 ;
        RECT 4.400 0.800 4.800 1.200 ;
      LAYER metal2 ;
        RECT 0.800 0.600 5.600 1.400 ;
      LAYER via2 ;
        RECT 1.600 0.800 2.000 1.200 ;
        RECT 3.000 0.800 3.400 1.200 ;
        RECT 4.400 0.800 4.800 1.200 ;
      LAYER metal3 ;
        RECT 0.800 0.400 5.600 1.600 ;
      LAYER via3 ;
        RECT 1.400 0.800 1.800 1.200 ;
        RECT 3.000 0.800 3.400 1.200 ;
        RECT 4.600 0.800 5.000 1.200 ;
      LAYER metal4 ;
        RECT 0.800 0.000 5.600 24.000 ;
    END
  END vdd
  PIN sum
    PORT
      LAYER metal1 ;
        RECT 14.000 14.300 14.800 19.800 ;
        RECT 17.200 14.300 18.000 14.400 ;
        RECT 14.000 13.700 18.000 14.300 ;
        RECT 14.000 12.400 14.800 13.700 ;
        RECT 17.200 13.600 18.000 13.700 ;
        RECT 14.200 10.200 14.800 12.400 ;
        RECT 14.000 2.200 14.800 10.200 ;
      LAYER via1 ;
        RECT 17.400 13.800 17.800 14.200 ;
      LAYER metal2 ;
        RECT 17.200 13.600 18.000 14.400 ;
        RECT 17.300 12.400 17.900 13.600 ;
        RECT 17.200 11.600 18.000 12.400 ;
      LAYER via2 ;
        RECT 17.400 11.800 17.800 12.200 ;
      LAYER metal3 ;
        RECT 17.200 11.600 18.000 12.400 ;
    END
  END sum
  PIN cout
    PORT
      LAYER metal1 ;
        RECT 1.200 14.300 2.000 14.400 ;
        RECT 6.000 14.300 6.800 19.800 ;
        RECT 1.200 13.700 6.800 14.300 ;
        RECT 1.200 13.600 2.000 13.700 ;
        RECT 6.000 12.400 6.800 13.700 ;
        RECT 6.000 10.200 6.600 12.400 ;
        RECT 6.000 2.200 6.800 10.200 ;
      LAYER via1 ;
        RECT 1.400 13.800 1.800 14.200 ;
      LAYER metal2 ;
        RECT 1.200 13.600 2.000 14.400 ;
        RECT 1.300 12.400 1.900 13.600 ;
        RECT 1.200 11.600 2.000 12.400 ;
      LAYER via2 ;
        RECT 1.400 11.800 1.800 12.200 ;
      LAYER metal3 ;
        RECT 1.200 12.300 2.000 12.400 ;
        RECT -1.900 11.700 2.000 12.300 ;
        RECT 1.200 11.600 2.000 11.700 ;
    END
  END cout
  OBS
      LAYER metal1 ;
        RECT 0.400 20.400 15.600 21.600 ;
        RECT 7.600 15.800 8.400 20.400 ;
        RECT 9.200 15.200 10.000 19.800 ;
        RECT 7.800 14.600 10.000 15.200 ;
        RECT 10.800 15.200 11.600 19.800 ;
        RECT 12.400 15.800 13.200 20.400 ;
        RECT 10.800 14.600 13.000 15.200 ;
        RECT 7.800 11.600 8.400 14.600 ;
        RECT 9.200 12.300 10.000 13.200 ;
        RECT 10.800 12.300 11.600 13.200 ;
        RECT 9.200 11.700 11.600 12.300 ;
        RECT 9.200 11.600 10.000 11.700 ;
        RECT 10.800 11.600 11.600 11.700 ;
        RECT 12.400 11.600 13.000 14.600 ;
        RECT 7.200 10.800 8.400 11.600 ;
        RECT 7.800 10.200 8.400 10.800 ;
        RECT 12.400 10.800 13.600 11.600 ;
        RECT 12.400 10.200 13.000 10.800 ;
        RECT 7.800 9.600 10.000 10.200 ;
        RECT 9.200 2.200 10.000 9.600 ;
        RECT 10.800 9.600 13.000 10.200 ;
        RECT 10.800 2.200 11.600 9.600 ;
      LAYER via1 ;
        RECT 7.800 16.000 8.200 16.400 ;
        RECT 9.400 11.800 9.800 12.200 ;
      LAYER metal2 ;
        RECT 7.600 16.300 8.400 16.600 ;
        RECT 7.600 15.800 9.900 16.300 ;
        RECT 7.700 15.700 9.900 15.800 ;
        RECT 9.300 12.400 9.900 15.700 ;
        RECT 9.200 11.600 10.000 12.400 ;
  END
END full_adder
END LIBRARY

