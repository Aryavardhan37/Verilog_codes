magic
tech scmos
timestamp 1706514480
<< metal1 >>
rect 200 103 202 107
rect 206 103 209 107
rect 213 103 216 107
rect 62 71 65 81
rect 270 72 273 81
rect 62 68 89 71
rect 158 68 169 71
rect 210 68 233 71
rect 86 62 89 68
rect 94 58 102 61
rect 126 58 137 61
rect 198 61 202 64
rect 198 58 206 61
rect 64 3 66 7
rect 70 3 73 7
rect 77 3 80 7
<< m2contact >>
rect 202 103 206 107
rect 209 103 213 107
rect 110 88 114 92
rect 262 88 266 92
rect 30 78 34 82
rect 6 68 10 72
rect 54 68 58 72
rect 142 78 146 82
rect 150 78 154 82
rect 182 68 186 72
rect 206 68 210 72
rect 238 68 242 72
rect 246 68 250 72
rect 270 68 274 72
rect 22 58 26 62
rect 46 58 50 62
rect 86 58 90 62
rect 102 58 106 62
rect 174 58 178 62
rect 190 58 194 62
rect 206 58 210 62
rect 222 58 226 62
rect 254 58 258 62
rect 102 48 106 52
rect 66 3 70 7
rect 73 3 77 7
<< metal2 >>
rect 94 102 97 131
rect 110 92 113 98
rect 150 92 153 131
rect 30 82 33 88
rect 150 82 153 88
rect 138 78 142 81
rect 50 68 54 71
rect 6 62 9 68
rect 22 62 25 68
rect 86 62 89 68
rect 50 58 54 61
rect 98 58 102 61
rect 134 52 137 78
rect 174 62 177 131
rect 200 103 202 107
rect 206 103 209 107
rect 213 103 216 107
rect 266 88 270 91
rect 182 72 185 78
rect 190 62 193 78
rect 206 72 209 88
rect 246 72 249 78
rect 270 72 273 78
rect 234 68 238 71
rect 218 58 222 61
rect 206 52 209 58
rect 254 52 257 58
rect 106 48 110 51
rect 64 3 66 7
rect 70 3 73 7
rect 77 3 80 7
<< m3contact >>
rect 94 98 98 102
rect 110 98 114 102
rect 30 88 34 92
rect 150 88 154 92
rect 134 78 138 82
rect 22 68 26 72
rect 46 68 50 72
rect 86 68 90 72
rect 6 58 10 62
rect 54 58 58 62
rect 94 58 98 62
rect 202 103 206 107
rect 209 103 213 107
rect 206 88 210 92
rect 270 88 274 92
rect 182 78 186 82
rect 190 78 194 82
rect 246 78 250 82
rect 270 78 274 82
rect 230 68 234 72
rect 174 58 178 62
rect 214 58 218 62
rect 254 58 258 62
rect 110 48 114 52
rect 134 48 138 52
rect 206 48 210 52
rect 254 48 258 52
rect 66 3 70 7
rect 73 3 77 7
<< metal3 >>
rect 200 103 202 107
rect 206 103 209 107
rect 214 103 216 107
rect 98 98 110 101
rect 154 88 206 91
rect 214 88 270 91
rect 30 81 33 88
rect -26 78 33 81
rect 138 78 182 81
rect 214 81 217 88
rect 194 78 217 81
rect 250 78 270 81
rect 274 78 305 81
rect 26 68 46 71
rect 90 68 230 71
rect -26 58 6 61
rect 58 58 94 61
rect 178 58 214 61
rect 258 58 305 61
rect 114 48 134 51
rect 210 48 254 51
rect 64 3 66 7
rect 70 3 73 7
rect 78 3 80 7
<< m4contact >>
rect 202 103 206 107
rect 210 103 213 107
rect 213 103 214 107
rect 66 3 70 7
rect 74 3 77 7
rect 77 3 78 7
<< metal4 >>
rect 200 103 202 107
rect 206 103 209 107
rect 214 103 216 107
rect 64 3 66 7
rect 70 3 73 7
rect 78 3 80 7
<< m5contact >>
rect 202 103 206 107
rect 209 103 210 107
rect 210 103 213 107
rect 66 3 70 7
rect 73 3 74 7
rect 74 3 77 7
<< metal5 >>
rect 206 103 209 107
rect 205 102 210 103
rect 215 102 216 107
rect 70 3 73 7
rect 69 2 74 3
rect 79 2 80 7
<< m6contact >>
rect 200 103 202 107
rect 202 103 205 107
rect 210 103 213 107
rect 213 103 215 107
rect 200 102 205 103
rect 210 102 215 103
rect 64 3 66 7
rect 66 3 69 7
rect 74 3 77 7
rect 77 3 79 7
rect 64 2 69 3
rect 74 2 79 3
<< metal6 >>
rect 64 7 80 130
rect 69 2 74 7
rect 79 2 80 7
rect 64 0 80 2
rect 200 107 216 130
rect 205 102 210 107
rect 215 102 216 107
rect 200 0 216 102
use BUFX2  BUFX2_2
timestamp 1706514480
transform -1 0 28 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_1
timestamp 1706514480
transform -1 0 52 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_3
timestamp 1706514480
transform -1 0 68 0 -1 105
box -2 -3 18 103
use FILL  FILL_0_0_0
timestamp 1706514480
transform 1 0 68 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1706514480
transform 1 0 76 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_1
timestamp 1706514480
transform 1 0 84 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_3
timestamp 1706514480
transform -1 0 132 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_2
timestamp 1706514480
transform -1 0 148 0 -1 105
box -2 -3 18 103
use INVX1  INVX1_4
timestamp 1706514480
transform 1 0 148 0 -1 105
box -2 -3 18 103
use OAI22X1  OAI22X1_1
timestamp 1706514480
transform 1 0 164 0 -1 105
box -2 -3 42 103
use FILL  FILL_0_1_0
timestamp 1706514480
transform 1 0 204 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1706514480
transform 1 0 212 0 -1 105
box -2 -3 10 103
use AOI22X1  AOI22X1_1
timestamp 1706514480
transform 1 0 220 0 -1 105
box -2 -3 42 103
use INVX1  INVX1_1
timestamp 1706514480
transform -1 0 276 0 -1 105
box -2 -3 18 103
<< labels >>
flabel metal6 s 64 0 80 8 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 200 0 216 8 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 176 130 176 130 3 FreeSans 24 90 0 0 x1
port 2 nsew
flabel metal3 s 304 80 304 80 3 FreeSans 24 270 0 0 x2
port 3 nsew
flabel metal2 s 152 130 152 130 3 FreeSans 24 90 0 0 x3
port 4 nsew
flabel metal3 s 304 60 304 60 3 FreeSans 24 270 0 0 x4
port 5 nsew
flabel metal3 s -24 60 -24 60 7 FreeSans 24 270 0 0 g
port 6 nsew
flabel metal2 s 96 130 96 130 3 FreeSans 24 90 0 0 h
port 7 nsew
flabel metal3 s -24 80 -24 80 7 FreeSans 24 270 0 0 f
port 8 nsew
<< end >>
