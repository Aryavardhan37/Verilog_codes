VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO down_counter_3bit
  CLASS BLOCK ;
  FOREIGN down_counter_3bit ;
  ORIGIN 1.900 4.000 ;
  SIZE 96.600 BY 48.300 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 0.400 40.400 92.400 41.600 ;
        RECT 2.800 33.000 3.600 40.400 ;
        RECT 7.800 39.800 8.600 40.400 ;
        RECT 7.600 33.200 8.600 39.800 ;
        RECT 13.800 33.200 14.800 40.400 ;
        RECT 22.000 35.800 22.800 40.400 ;
        RECT 25.200 35.800 26.000 40.400 ;
        RECT 28.400 35.800 29.200 40.400 ;
        RECT 31.600 35.800 32.400 40.400 ;
        RECT 39.600 35.800 40.400 40.400 ;
        RECT 42.800 35.800 43.600 40.400 ;
        RECT 49.200 35.800 50.000 40.400 ;
        RECT 52.400 35.800 53.200 40.400 ;
        RECT 55.600 35.800 56.400 40.400 ;
        RECT 58.800 35.800 59.600 40.400 ;
        RECT 49.000 31.800 49.800 32.000 ;
        RECT 52.400 31.800 53.200 32.400 ;
        RECT 60.400 31.800 61.200 40.400 ;
        RECT 64.600 35.800 65.400 40.400 ;
        RECT 71.600 35.800 72.400 40.400 ;
        RECT 74.800 35.800 75.600 40.400 ;
        RECT 78.000 36.200 78.800 40.400 ;
        RECT 81.200 35.800 82.000 40.400 ;
        RECT 84.400 35.800 85.200 40.400 ;
        RECT 87.600 33.000 88.400 40.400 ;
        RECT 26.200 31.200 53.200 31.800 ;
        RECT 26.200 31.000 27.000 31.200 ;
        RECT 5.400 10.800 6.200 11.000 ;
        RECT 73.800 10.800 74.600 11.000 ;
        RECT 5.400 10.200 32.400 10.800 ;
        RECT 47.600 10.200 74.600 10.800 ;
        RECT 28.200 10.000 29.200 10.200 ;
        RECT 31.600 9.600 32.400 10.200 ;
        RECT 1.200 1.600 2.000 6.200 ;
        RECT 4.400 1.600 5.200 6.200 ;
        RECT 7.600 1.600 8.400 6.200 ;
        RECT 10.800 1.600 11.600 6.200 ;
        RECT 18.800 1.600 19.600 6.200 ;
        RECT 22.000 1.600 22.800 6.200 ;
        RECT 28.400 1.600 29.200 6.200 ;
        RECT 31.600 1.600 32.400 6.200 ;
        RECT 34.800 1.600 35.600 6.200 ;
        RECT 42.800 1.600 43.600 10.200 ;
        RECT 47.600 9.600 48.400 10.200 ;
        RECT 51.000 10.000 51.800 10.200 ;
        RECT 44.400 1.600 45.200 6.200 ;
        RECT 47.600 1.600 48.400 6.200 ;
        RECT 50.800 1.600 51.600 6.200 ;
        RECT 57.200 1.600 58.000 6.200 ;
        RECT 60.400 1.600 61.200 6.200 ;
        RECT 68.400 1.600 69.200 6.200 ;
        RECT 71.600 1.600 72.400 6.200 ;
        RECT 74.800 1.600 75.600 6.200 ;
        RECT 78.000 1.600 78.800 6.200 ;
        RECT 86.000 1.600 86.800 6.200 ;
        RECT 89.200 1.600 90.000 9.000 ;
        RECT 0.400 0.400 92.400 1.600 ;
      LAYER via1 ;
        RECT 27.000 40.600 27.800 41.400 ;
        RECT 28.400 40.600 29.200 41.400 ;
        RECT 29.800 40.600 30.600 41.400 ;
        RECT 52.400 37.600 53.200 38.400 ;
        RECT 52.400 31.600 53.200 32.400 ;
        RECT 28.400 10.000 29.200 10.800 ;
        RECT 28.400 3.600 29.200 4.400 ;
        RECT 47.600 3.600 48.400 4.400 ;
        RECT 27.000 0.600 27.800 1.400 ;
        RECT 28.400 0.600 29.200 1.400 ;
        RECT 29.800 0.600 30.600 1.400 ;
      LAYER metal2 ;
        RECT 26.400 40.600 31.200 41.400 ;
        RECT 52.400 37.600 53.200 38.400 ;
        RECT 52.500 32.400 53.100 37.600 ;
        RECT 52.400 31.600 53.200 32.400 ;
        RECT 28.400 10.000 29.200 10.800 ;
        RECT 28.500 4.400 29.100 10.000 ;
        RECT 47.600 9.600 48.400 10.400 ;
        RECT 47.700 4.400 48.300 9.600 ;
        RECT 28.400 3.600 29.200 4.400 ;
        RECT 47.600 3.600 48.400 4.400 ;
        RECT 26.400 0.600 31.200 1.400 ;
      LAYER via2 ;
        RECT 27.000 40.600 27.800 41.400 ;
        RECT 28.400 40.600 29.200 41.400 ;
        RECT 29.800 40.600 30.600 41.400 ;
        RECT 27.000 0.600 27.800 1.400 ;
        RECT 28.400 0.600 29.200 1.400 ;
        RECT 29.800 0.600 30.600 1.400 ;
      LAYER metal3 ;
        RECT 26.400 40.400 31.200 41.600 ;
        RECT 26.400 0.400 31.200 1.600 ;
      LAYER via3 ;
        RECT 26.800 40.600 27.600 41.400 ;
        RECT 28.400 40.600 29.200 41.400 ;
        RECT 30.000 40.600 30.800 41.400 ;
        RECT 26.800 0.600 27.600 1.400 ;
        RECT 28.400 0.600 29.200 1.400 ;
        RECT 30.000 0.600 30.800 1.400 ;
      LAYER metal4 ;
        RECT 26.400 -4.000 31.200 44.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 2.800 21.600 3.600 26.200 ;
        RECT 7.600 22.200 8.600 25.600 ;
        RECT 7.800 21.600 8.600 22.200 ;
        RECT 13.800 21.600 14.800 25.600 ;
        RECT 22.000 21.600 22.800 24.200 ;
        RECT 28.400 21.600 29.200 26.200 ;
        RECT 39.600 21.600 40.400 24.200 ;
        RECT 42.800 21.600 43.600 24.200 ;
        RECT 52.400 21.600 53.200 26.200 ;
        RECT 58.800 21.600 59.600 24.200 ;
        RECT 62.000 21.600 62.800 25.400 ;
        RECT 71.600 21.600 72.400 26.200 ;
        RECT 81.200 21.600 82.000 28.200 ;
        RECT 84.400 21.600 85.200 24.200 ;
        RECT 87.600 21.600 88.400 26.200 ;
        RECT 0.400 20.400 92.400 21.600 ;
        RECT 1.200 17.800 2.000 20.400 ;
        RECT 7.600 15.800 8.400 20.400 ;
        RECT 18.800 17.800 19.600 20.400 ;
        RECT 22.000 17.800 22.800 20.400 ;
        RECT 31.600 15.800 32.400 20.400 ;
        RECT 42.800 15.800 43.600 20.400 ;
        RECT 47.600 15.800 48.400 20.400 ;
        RECT 57.200 17.800 58.000 20.400 ;
        RECT 60.400 17.800 61.200 20.400 ;
        RECT 71.600 15.800 72.400 20.400 ;
        RECT 78.000 17.800 78.800 20.400 ;
        RECT 86.000 17.800 86.800 20.400 ;
        RECT 89.200 15.800 90.000 20.400 ;
      LAYER via1 ;
        RECT 73.400 20.600 74.200 21.400 ;
        RECT 74.800 20.600 75.600 21.400 ;
        RECT 76.200 20.600 77.000 21.400 ;
      LAYER metal2 ;
        RECT 72.800 20.600 77.600 21.400 ;
      LAYER via2 ;
        RECT 73.400 20.600 74.200 21.400 ;
        RECT 74.800 20.600 75.600 21.400 ;
        RECT 76.200 20.600 77.000 21.400 ;
      LAYER metal3 ;
        RECT 72.800 20.400 77.600 21.600 ;
      LAYER via3 ;
        RECT 73.200 20.600 74.000 21.400 ;
        RECT 74.800 20.600 75.600 21.400 ;
        RECT 76.400 20.600 77.200 21.400 ;
      LAYER metal4 ;
        RECT 72.800 -4.000 77.600 44.000 ;
    END
  END gnd
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 38.800 25.600 40.400 26.400 ;
        RECT 18.000 15.600 19.600 16.400 ;
        RECT 60.400 15.600 62.000 16.400 ;
      LAYER via1 ;
        RECT 39.600 25.600 40.400 26.400 ;
        RECT 18.800 15.600 19.600 16.400 ;
      LAYER metal2 ;
        RECT 34.900 40.400 35.500 44.300 ;
        RECT 34.800 39.600 35.600 40.400 ;
        RECT 39.600 39.600 40.400 40.400 ;
        RECT 39.700 26.400 40.300 39.600 ;
        RECT 39.600 25.600 40.400 26.400 ;
        RECT 39.700 16.400 40.300 25.600 ;
        RECT 18.800 15.600 19.600 16.400 ;
        RECT 39.600 15.600 40.400 16.400 ;
        RECT 60.400 15.600 61.200 16.400 ;
      LAYER metal3 ;
        RECT 34.800 40.300 35.600 40.400 ;
        RECT 39.600 40.300 40.400 40.400 ;
        RECT 34.800 39.700 40.400 40.300 ;
        RECT 34.800 39.600 35.600 39.700 ;
        RECT 39.600 39.600 40.400 39.700 ;
        RECT 18.800 16.300 19.600 16.400 ;
        RECT 39.600 16.300 40.400 16.400 ;
        RECT 60.400 16.300 61.200 16.400 ;
        RECT 18.800 15.700 61.200 16.300 ;
        RECT 18.800 15.600 19.600 15.700 ;
        RECT 39.600 15.600 40.400 15.700 ;
        RECT 60.400 15.600 61.200 15.700 ;
    END
  END clk
  PIN rst
    PORT
      LAYER metal1 ;
        RECT 42.800 13.600 43.600 15.200 ;
      LAYER metal2 ;
        RECT 42.800 13.600 43.600 14.400 ;
        RECT 42.900 -1.700 43.500 13.600 ;
        RECT 41.300 -2.300 43.500 -1.700 ;
    END
  END rst
  PIN count[0]
    PORT
      LAYER metal1 ;
        RECT 1.200 31.800 2.000 39.800 ;
        RECT 1.200 29.600 1.800 31.800 ;
        RECT 1.200 22.200 2.000 29.600 ;
      LAYER via1 ;
        RECT 1.200 27.600 2.000 28.400 ;
      LAYER metal2 ;
        RECT 1.200 29.600 2.000 30.400 ;
        RECT 1.300 28.400 1.900 29.600 ;
        RECT 1.200 27.600 2.000 28.400 ;
      LAYER metal3 ;
        RECT 1.200 30.300 2.000 30.400 ;
        RECT -1.900 29.700 2.000 30.300 ;
        RECT 1.200 29.600 2.000 29.700 ;
    END
  END count[0]
  PIN count[1]
    PORT
      LAYER metal1 ;
        RECT 89.200 31.800 90.000 39.800 ;
        RECT 89.400 29.600 90.000 31.800 ;
        RECT 89.200 28.300 90.000 29.600 ;
        RECT 90.800 28.300 91.600 28.400 ;
        RECT 89.200 27.700 91.600 28.300 ;
        RECT 89.200 22.200 90.000 27.700 ;
        RECT 90.800 27.600 91.600 27.700 ;
      LAYER metal2 ;
        RECT 90.800 29.600 91.600 30.400 ;
        RECT 90.900 28.400 91.500 29.600 ;
        RECT 90.800 27.600 91.600 28.400 ;
      LAYER metal3 ;
        RECT 90.800 30.300 91.600 30.400 ;
        RECT 90.800 29.700 94.700 30.300 ;
        RECT 90.800 29.600 91.600 29.700 ;
    END
  END count[1]
  PIN count[2]
    PORT
      LAYER metal1 ;
        RECT 90.800 12.400 91.600 19.800 ;
        RECT 91.000 10.200 91.600 12.400 ;
        RECT 90.800 2.200 91.600 10.200 ;
      LAYER via1 ;
        RECT 90.800 7.600 91.600 8.400 ;
      LAYER metal2 ;
        RECT 90.800 9.600 91.600 10.400 ;
        RECT 90.900 8.400 91.500 9.600 ;
        RECT 90.800 7.600 91.600 8.400 ;
      LAYER metal3 ;
        RECT 90.800 10.300 91.600 10.400 ;
        RECT 90.800 9.700 94.700 10.300 ;
        RECT 90.800 9.600 91.600 9.700 ;
    END
  END count[2]
  OBS
      LAYER metal1 ;
        RECT 4.400 32.400 5.200 39.800 ;
        RECT 3.000 31.800 5.200 32.400 ;
        RECT 6.000 32.400 6.800 39.800 ;
        RECT 7.400 32.400 8.200 32.600 ;
        RECT 6.000 31.800 8.200 32.400 ;
        RECT 10.400 32.400 12.000 39.800 ;
        RECT 14.000 32.400 14.800 32.600 ;
        RECT 15.600 32.400 16.400 39.800 ;
        RECT 10.400 31.800 12.400 32.400 ;
        RECT 14.000 31.800 16.400 32.400 ;
        RECT 23.600 32.000 24.400 39.800 ;
        RECT 26.800 35.200 27.600 39.800 ;
        RECT 3.000 31.200 3.600 31.800 ;
        RECT 2.400 30.400 3.600 31.200 ;
        RECT 7.600 31.200 8.200 31.800 ;
        RECT 7.600 30.600 11.000 31.200 ;
        RECT 10.200 30.400 11.000 30.600 ;
        RECT 11.800 30.400 12.400 31.800 ;
        RECT 23.400 31.200 24.400 32.000 ;
        RECT 25.000 34.600 27.600 35.200 ;
        RECT 25.000 33.000 25.600 34.600 ;
        RECT 30.000 34.400 30.800 39.800 ;
        RECT 33.200 37.000 34.000 39.800 ;
        RECT 34.800 37.000 35.600 39.800 ;
        RECT 36.400 37.000 37.200 39.800 ;
        RECT 31.400 34.400 35.600 35.200 ;
        RECT 28.200 33.600 30.800 34.400 ;
        RECT 38.000 33.600 38.800 39.800 ;
        RECT 41.200 35.000 42.000 39.800 ;
        RECT 44.400 35.000 45.200 39.800 ;
        RECT 46.000 37.000 46.800 39.800 ;
        RECT 47.600 37.000 48.400 39.800 ;
        RECT 50.800 35.200 51.600 39.800 ;
        RECT 54.000 36.400 54.800 39.800 ;
        RECT 54.000 35.800 55.000 36.400 ;
        RECT 54.400 35.200 55.000 35.800 ;
        RECT 49.600 34.400 53.800 35.200 ;
        RECT 54.400 34.600 56.400 35.200 ;
        RECT 41.200 33.600 43.800 34.400 ;
        RECT 44.400 33.800 50.200 34.400 ;
        RECT 53.200 34.000 53.800 34.400 ;
        RECT 33.200 33.000 34.000 33.200 ;
        RECT 25.000 32.400 34.000 33.000 ;
        RECT 36.400 33.000 37.200 33.200 ;
        RECT 44.400 33.000 45.000 33.800 ;
        RECT 50.800 33.200 52.200 33.800 ;
        RECT 53.200 33.200 54.800 34.000 ;
        RECT 36.400 32.400 45.000 33.000 ;
        RECT 46.000 33.000 52.200 33.200 ;
        RECT 46.000 32.600 51.400 33.000 ;
        RECT 46.000 32.400 46.800 32.600 ;
        RECT 3.000 27.400 3.600 30.400 ;
        RECT 4.400 30.300 5.200 30.400 ;
        RECT 4.400 29.700 6.700 30.300 ;
        RECT 4.400 28.800 5.200 29.700 ;
        RECT 6.100 28.400 6.700 29.700 ;
        RECT 8.000 29.800 8.800 30.000 ;
        RECT 11.800 29.800 13.200 30.400 ;
        RECT 8.000 29.200 10.600 29.800 ;
        RECT 10.000 28.600 10.600 29.200 ;
        RECT 11.400 29.600 13.200 29.800 ;
        RECT 11.400 29.200 12.400 29.600 ;
        RECT 6.000 28.200 7.600 28.400 ;
        RECT 6.000 27.600 9.400 28.200 ;
        RECT 10.000 27.800 10.800 28.600 ;
        RECT 3.000 26.800 5.200 27.400 ;
        RECT 8.800 27.200 9.400 27.600 ;
        RECT 7.400 26.800 8.200 27.000 ;
        RECT 4.400 22.200 5.200 26.800 ;
        RECT 6.000 26.200 8.200 26.800 ;
        RECT 8.800 26.600 10.800 27.200 ;
        RECT 9.200 26.400 10.800 26.600 ;
        RECT 6.000 22.200 6.800 26.200 ;
        RECT 11.400 25.800 12.000 29.200 ;
        RECT 12.800 27.600 13.600 28.400 ;
        RECT 14.800 28.300 16.400 28.400 ;
        RECT 22.000 28.300 22.800 28.400 ;
        RECT 14.800 27.700 22.800 28.300 ;
        RECT 14.800 27.600 16.400 27.700 ;
        RECT 22.000 27.600 22.800 27.700 ;
        RECT 12.800 27.200 13.400 27.600 ;
        RECT 12.600 26.400 13.400 27.200 ;
        RECT 14.000 26.800 14.800 27.000 ;
        RECT 23.400 26.800 24.200 31.200 ;
        RECT 25.000 30.600 25.600 32.400 ;
        RECT 24.800 30.000 25.600 30.600 ;
        RECT 31.600 30.000 55.000 30.600 ;
        RECT 24.800 28.000 25.400 30.000 ;
        RECT 31.600 29.400 32.400 30.000 ;
        RECT 49.200 29.600 50.000 30.000 ;
        RECT 54.200 29.800 55.000 30.000 ;
        RECT 26.000 28.600 29.800 29.400 ;
        RECT 24.800 27.400 26.000 28.000 ;
        RECT 14.000 26.200 16.400 26.800 ;
        RECT 10.400 24.400 12.000 25.800 ;
        RECT 10.400 23.600 13.200 24.400 ;
        RECT 10.400 22.200 12.000 23.600 ;
        RECT 15.600 22.200 16.400 26.200 ;
        RECT 23.400 26.000 24.400 26.800 ;
        RECT 23.600 22.200 24.400 26.000 ;
        RECT 25.200 22.200 26.000 27.400 ;
        RECT 29.000 27.400 29.800 28.600 ;
        RECT 29.000 26.800 30.800 27.400 ;
        RECT 30.000 26.200 30.800 26.800 ;
        RECT 34.800 26.400 35.600 29.200 ;
        RECT 38.000 28.600 41.200 29.400 ;
        RECT 45.000 28.600 47.000 29.400 ;
        RECT 55.600 29.000 56.400 34.600 ;
        RECT 37.600 27.800 38.400 28.000 ;
        RECT 37.600 27.200 42.000 27.800 ;
        RECT 41.200 27.000 42.000 27.200 ;
        RECT 42.800 26.800 43.600 28.400 ;
        RECT 30.000 25.400 32.400 26.200 ;
        RECT 34.800 25.600 35.800 26.400 ;
        RECT 41.200 26.200 42.000 26.400 ;
        RECT 45.000 26.200 45.800 28.600 ;
        RECT 47.600 28.200 56.400 29.000 ;
        RECT 51.000 26.800 54.000 27.600 ;
        RECT 51.000 26.200 51.800 26.800 ;
        RECT 41.200 25.600 45.800 26.200 ;
        RECT 31.600 22.200 32.400 25.400 ;
        RECT 49.200 25.400 51.800 26.200 ;
        RECT 33.200 22.200 34.000 25.000 ;
        RECT 34.800 22.200 35.600 25.000 ;
        RECT 36.400 22.200 37.200 25.000 ;
        RECT 38.000 22.200 38.800 25.000 ;
        RECT 41.200 22.200 42.000 25.000 ;
        RECT 44.400 22.200 45.200 25.000 ;
        RECT 46.000 22.200 46.800 25.000 ;
        RECT 47.600 22.200 48.400 25.000 ;
        RECT 49.200 22.200 50.000 25.400 ;
        RECT 55.600 22.200 56.400 28.200 ;
        RECT 57.200 22.200 58.000 39.800 ;
        RECT 63.000 32.400 63.800 39.800 ;
        RECT 64.400 33.600 65.200 34.400 ;
        RECT 64.600 32.400 65.200 33.600 ;
        RECT 63.000 31.800 64.000 32.400 ;
        RECT 64.600 32.300 66.000 32.400 ;
        RECT 68.400 32.300 69.200 32.400 ;
        RECT 64.600 31.800 69.200 32.300 ;
        RECT 62.000 28.800 62.800 30.400 ;
        RECT 63.400 28.400 64.000 31.800 ;
        RECT 65.200 31.700 69.200 31.800 ;
        RECT 65.200 31.600 66.000 31.700 ;
        RECT 68.400 31.600 69.200 31.700 ;
        RECT 60.400 28.300 61.200 28.400 ;
        RECT 58.900 28.200 61.200 28.300 ;
        RECT 63.400 28.300 66.000 28.400 ;
        RECT 71.600 28.300 72.400 28.400 ;
        RECT 58.900 27.700 62.000 28.200 ;
        RECT 58.900 26.400 59.500 27.700 ;
        RECT 60.400 27.600 62.000 27.700 ;
        RECT 63.400 27.700 72.400 28.300 ;
        RECT 63.400 27.600 66.000 27.700 ;
        RECT 61.200 27.200 62.000 27.600 ;
        RECT 58.800 24.800 59.600 26.400 ;
        RECT 60.600 26.200 64.200 26.600 ;
        RECT 65.200 26.200 65.800 27.600 ;
        RECT 71.600 26.800 72.400 27.700 ;
        RECT 73.200 26.200 74.000 39.800 ;
        RECT 76.400 35.800 77.200 39.800 ;
        RECT 76.600 35.600 77.200 35.800 ;
        RECT 79.600 35.800 80.400 39.800 ;
        RECT 79.600 35.600 80.200 35.800 ;
        RECT 76.600 35.000 80.200 35.600 ;
        RECT 74.800 32.300 75.600 33.200 ;
        RECT 76.600 32.400 77.200 35.000 ;
        RECT 78.000 34.300 78.800 34.400 ;
        RECT 82.800 34.300 83.600 39.800 ;
        RECT 78.000 33.700 83.600 34.300 ;
        RECT 78.000 32.800 78.800 33.700 ;
        RECT 76.400 32.300 77.200 32.400 ;
        RECT 74.800 31.700 77.200 32.300 ;
        RECT 74.800 31.600 75.600 31.700 ;
        RECT 76.400 31.600 77.200 31.700 ;
        RECT 76.600 28.400 77.200 31.600 ;
        RECT 78.000 29.600 80.400 30.400 ;
        RECT 81.200 29.600 82.000 32.400 ;
        RECT 76.600 28.200 78.200 28.400 ;
        RECT 76.600 27.800 78.400 28.200 ;
        RECT 60.400 26.000 64.400 26.200 ;
        RECT 60.400 22.200 61.200 26.000 ;
        RECT 63.600 22.200 64.400 26.000 ;
        RECT 65.200 22.200 66.000 26.200 ;
        RECT 73.200 25.600 75.000 26.200 ;
        RECT 74.200 24.400 75.000 25.600 ;
        RECT 73.200 23.600 75.000 24.400 ;
        RECT 74.200 22.200 75.000 23.600 ;
        RECT 77.600 22.200 78.400 27.800 ;
        RECT 82.800 22.200 83.600 33.700 ;
        RECT 86.000 32.400 86.800 39.800 ;
        RECT 86.000 31.800 88.200 32.400 ;
        RECT 87.600 31.200 88.200 31.800 ;
        RECT 87.600 30.400 88.800 31.200 ;
        RECT 84.400 30.300 85.200 30.400 ;
        RECT 86.000 30.300 86.800 30.400 ;
        RECT 84.400 29.700 86.800 30.300 ;
        RECT 84.400 29.600 85.200 29.700 ;
        RECT 86.000 28.800 86.800 29.700 ;
        RECT 87.600 27.400 88.200 30.400 ;
        RECT 86.000 26.800 88.200 27.400 ;
        RECT 84.400 24.800 85.200 26.400 ;
        RECT 86.000 22.200 86.800 26.800 ;
        RECT 2.800 16.000 3.600 19.800 ;
        RECT 2.600 15.200 3.600 16.000 ;
        RECT 2.600 10.800 3.400 15.200 ;
        RECT 4.400 14.600 5.200 19.800 ;
        RECT 10.800 16.600 11.600 19.800 ;
        RECT 12.400 17.000 13.200 19.800 ;
        RECT 14.000 17.000 14.800 19.800 ;
        RECT 15.600 17.000 16.400 19.800 ;
        RECT 17.200 17.000 18.000 19.800 ;
        RECT 20.400 17.000 21.200 19.800 ;
        RECT 23.600 17.000 24.400 19.800 ;
        RECT 25.200 17.000 26.000 19.800 ;
        RECT 26.800 17.000 27.600 19.800 ;
        RECT 9.200 15.800 11.600 16.600 ;
        RECT 28.400 16.600 29.200 19.800 ;
        RECT 9.200 15.200 10.000 15.800 ;
        RECT 4.000 14.000 5.200 14.600 ;
        RECT 8.200 14.600 10.000 15.200 ;
        RECT 14.000 15.600 15.000 16.400 ;
        RECT 20.400 15.800 25.000 16.400 ;
        RECT 28.400 15.800 31.000 16.600 ;
        RECT 20.400 15.600 21.200 15.800 ;
        RECT 4.000 12.000 4.600 14.000 ;
        RECT 8.200 13.400 9.000 14.600 ;
        RECT 5.200 12.600 9.000 13.400 ;
        RECT 14.000 12.800 14.800 15.600 ;
        RECT 20.400 14.800 21.200 15.000 ;
        RECT 16.800 14.200 21.200 14.800 ;
        RECT 16.800 14.000 17.600 14.200 ;
        RECT 22.000 13.600 22.800 15.200 ;
        RECT 24.200 13.400 25.000 15.800 ;
        RECT 30.200 15.200 31.000 15.800 ;
        RECT 30.200 14.400 33.200 15.200 ;
        RECT 34.800 13.800 35.600 19.800 ;
        RECT 17.200 12.600 20.400 13.400 ;
        RECT 24.200 12.600 26.200 13.400 ;
        RECT 26.800 13.000 35.600 13.800 ;
        RECT 10.800 12.000 11.600 12.600 ;
        RECT 28.400 12.000 29.200 12.400 ;
        RECT 31.600 12.000 32.400 12.400 ;
        RECT 33.400 12.000 34.200 12.200 ;
        RECT 4.000 11.400 4.800 12.000 ;
        RECT 10.800 11.400 34.200 12.000 ;
        RECT 2.600 10.000 3.600 10.800 ;
        RECT 2.800 2.200 3.600 10.000 ;
        RECT 4.200 9.600 4.800 11.400 ;
        RECT 4.200 9.000 13.200 9.600 ;
        RECT 4.200 7.400 4.800 9.000 ;
        RECT 12.400 8.800 13.200 9.000 ;
        RECT 15.600 9.000 24.200 9.600 ;
        RECT 15.600 8.800 16.400 9.000 ;
        RECT 7.400 7.600 10.000 8.400 ;
        RECT 4.200 6.800 6.800 7.400 ;
        RECT 6.000 2.200 6.800 6.800 ;
        RECT 9.200 2.200 10.000 7.600 ;
        RECT 10.600 6.800 14.800 7.600 ;
        RECT 12.400 2.200 13.200 5.000 ;
        RECT 14.000 2.200 14.800 5.000 ;
        RECT 15.600 2.200 16.400 5.000 ;
        RECT 17.200 2.200 18.000 8.400 ;
        RECT 20.400 7.600 23.000 8.400 ;
        RECT 23.600 8.200 24.200 9.000 ;
        RECT 25.200 9.400 26.000 9.600 ;
        RECT 25.200 9.000 30.600 9.400 ;
        RECT 25.200 8.800 31.400 9.000 ;
        RECT 30.000 8.200 31.400 8.800 ;
        RECT 23.600 7.600 29.400 8.200 ;
        RECT 32.400 8.000 34.000 8.800 ;
        RECT 32.400 7.600 33.000 8.000 ;
        RECT 20.400 2.200 21.200 7.000 ;
        RECT 23.600 2.200 24.400 7.000 ;
        RECT 28.800 6.800 33.000 7.600 ;
        RECT 34.800 7.400 35.600 13.000 ;
        RECT 33.600 6.800 35.600 7.400 ;
        RECT 25.200 2.200 26.000 5.000 ;
        RECT 26.800 2.200 27.600 5.000 ;
        RECT 30.000 2.200 30.800 6.800 ;
        RECT 33.600 6.200 34.200 6.800 ;
        RECT 33.200 5.600 34.200 6.200 ;
        RECT 33.200 2.200 34.000 5.600 ;
        RECT 41.200 2.200 42.000 19.800 ;
        RECT 44.400 13.800 45.200 19.800 ;
        RECT 50.800 16.600 51.600 19.800 ;
        RECT 52.400 17.000 53.200 19.800 ;
        RECT 54.000 17.000 54.800 19.800 ;
        RECT 55.600 17.000 56.400 19.800 ;
        RECT 58.800 17.000 59.600 19.800 ;
        RECT 62.000 17.000 62.800 19.800 ;
        RECT 63.600 17.000 64.400 19.800 ;
        RECT 65.200 17.000 66.000 19.800 ;
        RECT 66.800 17.000 67.600 19.800 ;
        RECT 49.000 15.800 51.600 16.600 ;
        RECT 68.400 16.600 69.200 19.800 ;
        RECT 55.000 15.800 59.600 16.400 ;
        RECT 49.000 15.200 49.800 15.800 ;
        RECT 46.800 14.400 49.800 15.200 ;
        RECT 44.400 13.000 53.200 13.800 ;
        RECT 55.000 13.400 55.800 15.800 ;
        RECT 58.800 15.600 59.600 15.800 ;
        RECT 65.000 15.600 66.000 16.400 ;
        RECT 68.400 15.800 70.800 16.600 ;
        RECT 57.200 13.600 58.000 15.200 ;
        RECT 58.800 14.800 59.600 15.000 ;
        RECT 58.800 14.200 63.200 14.800 ;
        RECT 62.400 14.000 63.200 14.200 ;
        RECT 44.400 7.400 45.200 13.000 ;
        RECT 53.800 12.600 55.800 13.400 ;
        RECT 59.600 12.600 62.800 13.400 ;
        RECT 65.200 12.800 66.000 15.600 ;
        RECT 70.000 15.200 70.800 15.800 ;
        RECT 70.000 14.600 71.800 15.200 ;
        RECT 71.000 13.400 71.800 14.600 ;
        RECT 74.800 14.600 75.600 19.800 ;
        RECT 76.400 16.000 77.200 19.800 ;
        RECT 81.200 18.300 82.000 18.400 ;
        RECT 84.400 18.300 85.200 19.800 ;
        RECT 81.200 17.700 85.200 18.300 ;
        RECT 81.200 17.600 82.000 17.700 ;
        RECT 76.400 15.200 77.400 16.000 ;
        RECT 74.800 14.000 76.000 14.600 ;
        RECT 71.000 12.600 74.800 13.400 ;
        RECT 45.800 12.000 46.600 12.200 ;
        RECT 47.600 12.000 48.400 12.400 ;
        RECT 50.800 12.000 51.600 12.400 ;
        RECT 68.400 12.000 69.200 12.600 ;
        RECT 75.400 12.000 76.000 14.000 ;
        RECT 45.800 11.400 69.200 12.000 ;
        RECT 75.200 11.400 76.000 12.000 ;
        RECT 75.200 9.600 75.800 11.400 ;
        RECT 76.600 10.800 77.400 15.200 ;
        RECT 54.000 9.400 54.800 9.600 ;
        RECT 49.400 9.000 54.800 9.400 ;
        RECT 48.600 8.800 54.800 9.000 ;
        RECT 55.800 9.000 64.400 9.600 ;
        RECT 46.000 8.000 47.600 8.800 ;
        RECT 48.600 8.200 50.000 8.800 ;
        RECT 55.800 8.200 56.400 9.000 ;
        RECT 63.600 8.800 64.400 9.000 ;
        RECT 66.800 9.000 75.800 9.600 ;
        RECT 66.800 8.800 67.600 9.000 ;
        RECT 47.000 7.600 47.600 8.000 ;
        RECT 50.600 7.600 56.400 8.200 ;
        RECT 57.000 7.600 59.600 8.400 ;
        RECT 44.400 6.800 46.400 7.400 ;
        RECT 47.000 6.800 51.200 7.600 ;
        RECT 45.800 6.200 46.400 6.800 ;
        RECT 45.800 5.600 46.800 6.200 ;
        RECT 46.000 2.200 46.800 5.600 ;
        RECT 49.200 2.200 50.000 6.800 ;
        RECT 52.400 2.200 53.200 5.000 ;
        RECT 54.000 2.200 54.800 5.000 ;
        RECT 55.600 2.200 56.400 7.000 ;
        RECT 58.800 2.200 59.600 7.000 ;
        RECT 62.000 2.200 62.800 8.400 ;
        RECT 70.000 7.600 72.600 8.400 ;
        RECT 65.200 6.800 69.400 7.600 ;
        RECT 63.600 2.200 64.400 5.000 ;
        RECT 65.200 2.200 66.000 5.000 ;
        RECT 66.800 2.200 67.600 5.000 ;
        RECT 70.000 2.200 70.800 7.600 ;
        RECT 75.200 7.400 75.800 9.000 ;
        RECT 73.200 6.800 75.800 7.400 ;
        RECT 76.400 10.000 77.400 10.800 ;
        RECT 73.200 2.200 74.000 6.800 ;
        RECT 76.400 2.200 77.200 10.000 ;
        RECT 84.400 2.200 85.200 17.700 ;
        RECT 86.000 15.600 86.800 17.200 ;
        RECT 87.600 15.200 88.400 19.800 ;
        RECT 87.600 14.600 89.800 15.200 ;
        RECT 86.000 12.300 86.800 12.400 ;
        RECT 87.600 12.300 88.400 13.200 ;
        RECT 86.000 11.700 88.400 12.300 ;
        RECT 86.000 11.600 86.800 11.700 ;
        RECT 87.600 11.600 88.400 11.700 ;
        RECT 89.200 11.600 89.800 14.600 ;
        RECT 89.200 10.800 90.400 11.600 ;
        RECT 89.200 10.200 89.800 10.800 ;
        RECT 87.600 9.600 89.800 10.200 ;
        RECT 87.600 2.200 88.400 9.600 ;
      LAYER via1 ;
        RECT 7.400 31.800 8.200 32.600 ;
        RECT 34.800 34.400 35.600 35.200 ;
        RECT 38.000 35.000 38.800 35.800 ;
        RECT 33.200 32.400 34.000 33.200 ;
        RECT 7.400 26.200 8.200 27.000 ;
        RECT 31.600 29.600 32.400 30.400 ;
        RECT 12.400 23.600 13.200 24.400 ;
        RECT 23.600 25.600 24.400 26.400 ;
        RECT 42.800 27.600 43.600 28.400 ;
        RECT 33.200 24.200 34.000 25.000 ;
        RECT 34.800 24.200 35.600 25.000 ;
        RECT 36.400 24.200 37.200 25.000 ;
        RECT 38.000 24.200 38.800 25.000 ;
        RECT 41.200 24.200 42.000 25.000 ;
        RECT 44.400 24.200 45.200 25.000 ;
        RECT 46.000 24.200 46.800 25.000 ;
        RECT 47.600 24.200 48.400 25.000 ;
        RECT 62.000 29.600 62.800 30.400 ;
        RECT 57.200 27.600 58.000 28.400 ;
        RECT 58.800 25.600 59.600 26.400 ;
        RECT 84.400 25.600 85.200 26.400 ;
        RECT 2.800 17.600 3.600 18.400 ;
        RECT 20.400 14.200 21.200 15.000 ;
        RECT 31.600 11.600 32.400 12.400 ;
        RECT 14.000 6.800 14.800 7.600 ;
        RECT 17.200 6.200 18.000 7.000 ;
        RECT 12.400 4.200 13.200 5.000 ;
        RECT 14.000 4.200 14.800 5.000 ;
        RECT 15.600 4.200 16.400 5.000 ;
        RECT 20.400 6.200 21.200 7.000 ;
        RECT 23.600 6.200 24.400 7.000 ;
        RECT 41.200 11.600 42.000 12.400 ;
        RECT 25.200 4.200 26.000 5.000 ;
        RECT 26.800 4.200 27.600 5.000 ;
        RECT 52.400 13.000 53.200 13.800 ;
        RECT 62.000 12.600 62.800 13.400 ;
        RECT 47.600 11.600 48.400 12.400 ;
        RECT 76.600 11.600 77.400 12.400 ;
        RECT 54.000 8.800 54.800 9.600 ;
        RECT 58.800 7.600 59.600 8.400 ;
        RECT 55.600 6.200 56.400 7.000 ;
        RECT 52.400 4.200 53.200 5.000 ;
        RECT 54.000 4.200 54.800 5.000 ;
        RECT 58.800 6.200 59.600 7.000 ;
        RECT 62.000 6.200 62.800 7.000 ;
        RECT 63.600 4.200 64.400 5.000 ;
        RECT 65.200 4.200 66.000 5.000 ;
        RECT 66.800 4.200 67.600 5.000 ;
      LAYER metal2 ;
        RECT 7.400 31.800 8.200 32.600 ;
        RECT 14.000 31.800 14.800 32.600 ;
        RECT 2.800 29.600 3.600 30.400 ;
        RECT 2.900 18.400 3.500 29.600 ;
        RECT 7.400 27.000 8.000 31.800 ;
        RECT 10.000 28.400 10.800 28.600 ;
        RECT 14.200 28.400 14.800 31.800 ;
        RECT 22.000 29.600 22.800 30.400 ;
        RECT 31.600 29.600 32.400 30.400 ;
        RECT 22.100 28.400 22.700 29.600 ;
        RECT 10.000 27.800 14.800 28.400 ;
        RECT 9.200 27.000 10.000 27.200 ;
        RECT 12.600 27.000 13.400 27.200 ;
        RECT 14.200 27.000 14.800 27.800 ;
        RECT 22.000 27.600 22.800 28.400 ;
        RECT 7.400 26.200 8.200 27.000 ;
        RECT 9.200 26.400 13.400 27.000 ;
        RECT 12.400 25.600 13.200 26.400 ;
        RECT 14.000 26.200 14.800 27.000 ;
        RECT 23.600 25.600 24.400 26.400 ;
        RECT 12.400 23.600 13.200 24.400 ;
        RECT 22.000 23.600 22.800 24.400 ;
        RECT 2.800 17.600 3.600 18.400 ;
        RECT 12.400 4.200 13.200 17.800 ;
        RECT 14.000 4.200 14.800 17.800 ;
        RECT 15.600 4.200 16.400 17.800 ;
        RECT 17.200 6.200 18.000 17.800 ;
        RECT 20.400 6.200 21.200 17.800 ;
        RECT 22.100 14.400 22.700 23.600 ;
        RECT 22.000 13.600 22.800 14.400 ;
        RECT 23.600 6.200 24.400 17.800 ;
        RECT 25.200 4.200 26.000 17.800 ;
        RECT 26.800 4.200 27.600 17.800 ;
        RECT 31.700 12.400 32.300 29.600 ;
        RECT 33.200 24.200 34.000 37.800 ;
        RECT 34.800 24.200 35.600 37.800 ;
        RECT 36.400 24.200 37.200 37.800 ;
        RECT 38.000 24.200 38.800 35.800 ;
        RECT 41.200 24.200 42.000 35.800 ;
        RECT 42.800 27.600 43.600 28.400 ;
        RECT 44.400 24.200 45.200 35.800 ;
        RECT 46.000 24.200 46.800 37.800 ;
        RECT 47.600 24.200 48.400 37.800 ;
        RECT 68.400 31.600 69.200 32.400 ;
        RECT 62.000 29.600 62.800 30.400 ;
        RECT 57.200 27.600 58.000 28.400 ;
        RECT 58.800 25.600 59.600 26.400 ;
        RECT 57.200 23.600 58.000 24.400 ;
        RECT 31.600 11.600 32.400 12.400 ;
        RECT 41.200 11.600 42.000 12.400 ;
        RECT 47.600 11.600 48.400 12.400 ;
        RECT 52.400 4.200 53.200 17.800 ;
        RECT 54.000 4.200 54.800 17.800 ;
        RECT 55.600 6.200 56.400 17.800 ;
        RECT 57.300 14.400 57.900 23.600 ;
        RECT 57.200 13.600 58.000 14.400 ;
        RECT 58.800 6.200 59.600 17.800 ;
        RECT 62.000 6.200 62.800 17.800 ;
        RECT 63.600 4.200 64.400 17.800 ;
        RECT 65.200 4.200 66.000 17.800 ;
        RECT 66.800 4.200 67.600 17.800 ;
        RECT 68.500 12.400 69.100 31.600 ;
        RECT 78.000 29.600 78.800 30.400 ;
        RECT 81.200 29.600 82.000 30.400 ;
        RECT 84.400 29.600 85.200 30.400 ;
        RECT 78.100 28.400 78.700 29.600 ;
        RECT 78.000 27.600 78.800 28.400 ;
        RECT 73.200 23.600 74.000 24.400 ;
        RECT 81.300 18.400 81.900 29.600 ;
        RECT 84.500 26.400 85.100 29.600 ;
        RECT 84.400 25.600 85.200 26.400 ;
        RECT 81.200 17.600 82.000 18.400 ;
        RECT 86.000 15.600 86.800 16.400 ;
        RECT 86.100 12.400 86.700 15.600 ;
        RECT 68.400 11.600 69.200 12.400 ;
        RECT 76.400 11.600 77.400 12.400 ;
        RECT 86.000 11.600 86.800 12.400 ;
      LAYER via2 ;
        RECT 76.400 11.600 77.200 12.400 ;
      LAYER metal3 ;
        RECT 2.800 30.300 3.600 30.400 ;
        RECT 22.000 30.300 22.800 30.400 ;
        RECT 62.000 30.300 62.800 30.400 ;
        RECT 84.400 30.300 85.200 30.400 ;
        RECT 2.800 29.700 85.200 30.300 ;
        RECT 2.800 29.600 3.600 29.700 ;
        RECT 22.000 29.600 22.800 29.700 ;
        RECT 62.000 29.600 62.800 29.700 ;
        RECT 84.400 29.600 85.200 29.700 ;
        RECT 42.800 28.300 43.600 28.400 ;
        RECT 57.200 28.300 58.000 28.400 ;
        RECT 78.000 28.300 78.800 28.400 ;
        RECT 42.800 27.700 78.800 28.300 ;
        RECT 42.800 27.600 43.600 27.700 ;
        RECT 57.200 27.600 58.000 27.700 ;
        RECT 78.000 27.600 78.800 27.700 ;
        RECT 12.400 26.300 13.200 26.400 ;
        RECT 23.600 26.300 24.400 26.400 ;
        RECT 58.800 26.300 59.600 26.400 ;
        RECT 12.400 25.700 59.600 26.300 ;
        RECT 12.400 25.600 13.200 25.700 ;
        RECT 23.600 25.600 24.400 25.700 ;
        RECT 58.800 25.600 59.600 25.700 ;
        RECT 12.400 24.300 13.200 24.400 ;
        RECT 22.000 24.300 22.800 24.400 ;
        RECT 12.400 23.700 22.800 24.300 ;
        RECT 12.400 23.600 13.200 23.700 ;
        RECT 22.000 23.600 22.800 23.700 ;
        RECT 57.200 24.300 58.000 24.400 ;
        RECT 73.200 24.300 74.000 24.400 ;
        RECT 57.200 23.700 74.000 24.300 ;
        RECT 57.200 23.600 58.000 23.700 ;
        RECT 73.200 23.600 74.000 23.700 ;
        RECT 31.600 12.300 32.400 12.400 ;
        RECT 41.200 12.300 42.000 12.400 ;
        RECT 47.600 12.300 48.400 12.400 ;
        RECT 31.600 11.700 48.400 12.300 ;
        RECT 31.600 11.600 32.400 11.700 ;
        RECT 41.200 11.600 42.000 11.700 ;
        RECT 47.600 11.600 48.400 11.700 ;
        RECT 68.400 12.300 69.200 12.400 ;
        RECT 76.400 12.300 77.200 12.400 ;
        RECT 86.000 12.300 86.800 12.400 ;
        RECT 68.400 11.700 86.800 12.300 ;
        RECT 68.400 11.600 69.200 11.700 ;
        RECT 76.400 11.600 77.200 11.700 ;
        RECT 86.000 11.600 86.800 11.700 ;
  END
END down_counter_3bit
END LIBRARY

