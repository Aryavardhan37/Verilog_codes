module or_gate(a,b,y);
input a,b;
output y;
or(y,a,b);
endmodule