* NGSPICE file created from down_counter_3bit.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

.subckt down_counter_3bit vdd gnd clk rst count[0] count[1] count[2]
XFILL_0_0_0 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XFILL_0_0_2 gnd vdd FILL
XNAND3X1_1 INVX1_2/Y DFFSR_1/D INVX1_1/Y gnd NAND2X1_1/B vdd NAND3X1
XFILL_1_1_0 gnd vdd FILL
XFILL_1_1_1 gnd vdd FILL
XFILL_1_1_2 gnd vdd FILL
XOAI21X1_1 INVX1_3/A BUFX2_2/A BUFX2_3/A gnd NAND2X1_1/A vdd OAI21X1
XBUFX2_1 INVX1_3/A gnd count[0] vdd BUFX2
XBUFX2_2 BUFX2_2/A gnd count[1] vdd BUFX2
XINVX2_1 rst gnd DFFSR_1/R vdd INVX2
XBUFX2_3 BUFX2_3/A gnd count[2] vdd BUFX2
XFILL_0_1_0 gnd vdd FILL
XNAND2X1_1 NAND2X1_1/A NAND2X1_1/B gnd DFFSR_3/D vdd NAND2X1
XFILL_0_1_1 gnd vdd FILL
XFILL_0_1_2 gnd vdd FILL
XFILL_1_0_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XFILL_1_0_2 gnd vdd FILL
XDFFSR_1 INVX1_3/A clk DFFSR_1/R vdd DFFSR_1/D gnd vdd DFFSR
XDFFSR_3 BUFX2_3/A clk DFFSR_1/R vdd DFFSR_3/D gnd vdd DFFSR
XDFFSR_2 BUFX2_2/A clk DFFSR_1/R vdd DFFSR_2/D gnd vdd DFFSR
XFILL_2_1 gnd vdd FILL
XINVX1_1 BUFX2_2/A gnd INVX1_1/Y vdd INVX1
XXNOR2X1_1 INVX1_3/A BUFX2_2/A gnd DFFSR_2/D vdd XNOR2X1
XINVX1_2 BUFX2_3/A gnd INVX1_2/Y vdd INVX1
XINVX1_3 INVX1_3/A gnd DFFSR_1/D vdd INVX1
.ends

