module xnor_gate(a,b,y);
input a,b;
output y;
xnor(y,a,b);
endmodule