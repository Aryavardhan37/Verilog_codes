magic
tech scmos
timestamp 1697958199
<< metal1 >>
rect 96 103 98 107
rect 102 103 105 107
rect 109 103 112 107
rect 42 78 49 81
rect 14 68 30 71
rect 94 68 124 71
rect 62 58 73 61
rect 142 56 146 58
rect 126 38 134 41
rect 24 3 26 7
rect 30 3 33 7
rect 37 3 40 7
<< m2contact >>
rect 98 103 102 107
rect 105 103 109 107
rect 38 78 42 82
rect 6 68 10 72
rect 30 68 34 72
rect 86 66 90 70
rect 134 58 138 62
rect 142 58 146 62
rect 22 48 26 52
rect 134 38 138 42
rect 26 3 30 7
rect 33 3 37 7
<< metal2 >>
rect 96 103 98 107
rect 102 103 105 107
rect 109 103 112 107
rect 6 72 9 98
rect 34 78 38 81
rect 34 68 38 71
rect 82 66 86 69
rect 134 62 137 78
rect 22 52 25 58
rect 142 52 145 58
rect 138 38 142 41
rect 24 3 26 7
rect 30 3 33 7
rect 37 3 40 7
<< m3contact >>
rect 98 103 102 107
rect 105 103 109 107
rect 6 98 10 102
rect 30 78 34 82
rect 134 78 138 82
rect 38 68 42 72
rect 78 66 82 70
rect 22 58 26 62
rect 142 48 146 52
rect 142 38 146 42
rect 26 3 30 7
rect 33 3 37 7
<< metal3 >>
rect 96 103 98 107
rect 102 103 105 107
rect 110 103 112 107
rect -26 98 6 101
rect -26 78 30 81
rect 138 78 177 81
rect 42 70 81 71
rect 42 68 78 70
rect -26 58 22 61
rect 142 58 177 61
rect 142 52 145 58
rect 146 38 177 41
rect 24 3 26 7
rect 30 3 33 7
rect 38 3 40 7
<< m4contact >>
rect 98 103 102 107
rect 106 103 109 107
rect 109 103 110 107
rect 26 3 30 7
rect 34 3 37 7
rect 37 3 38 7
<< metal4 >>
rect 96 103 98 107
rect 102 103 105 107
rect 110 103 112 107
rect 24 3 26 7
rect 30 3 33 7
rect 38 3 40 7
<< m5contact >>
rect 98 103 102 107
rect 105 103 106 107
rect 106 103 109 107
rect 26 3 30 7
rect 33 3 34 7
rect 34 3 37 7
<< metal5 >>
rect 102 103 105 107
rect 101 102 106 103
rect 111 102 112 107
rect 30 3 33 7
rect 29 2 34 3
rect 39 2 40 7
<< m6contact >>
rect 96 103 98 107
rect 98 103 101 107
rect 106 103 109 107
rect 109 103 111 107
rect 96 102 101 103
rect 106 102 111 103
rect 24 3 26 7
rect 26 3 29 7
rect 34 3 37 7
rect 37 3 39 7
rect 24 2 29 3
rect 34 2 39 3
<< metal6 >>
rect 24 7 40 110
rect 29 2 34 7
rect 39 2 40 7
rect 24 0 40 2
rect 96 107 112 110
rect 101 102 106 107
rect 111 102 112 107
rect 96 0 112 102
use NAND3X1  NAND3X1_1
timestamp 1697958199
transform -1 0 148 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_1_1
timestamp 1697958199
transform -1 0 116 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_0
timestamp 1697958199
transform -1 0 108 0 -1 105
box -2 -3 10 103
use AND2X2  AND2X2_1
timestamp 1697958199
transform -1 0 100 0 -1 105
box -2 -3 34 103
use BUFX2  BUFX2_1
timestamp 1697958199
transform -1 0 68 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_0_1
timestamp 1697958199
transform -1 0 44 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_0
timestamp 1697958199
transform -1 0 36 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_1
timestamp 1697958199
transform 1 0 4 0 -1 105
box -2 -3 26 103
<< labels >>
flabel metal6 s 24 0 40 8 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 96 0 112 8 3 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal3 s -24 60 -24 60 7 FreeSans 24 270 0 0 A
port 2 nsew
flabel metal3 s -24 100 -24 100 7 FreeSans 24 270 0 0 B
port 3 nsew
flabel metal3 s 176 80 176 80 3 FreeSans 24 270 0 0 C
port 4 nsew
flabel metal3 s 176 60 176 60 3 FreeSans 24 270 0 0 D
port 5 nsew
flabel metal3 s 176 40 176 40 3 FreeSans 24 270 0 0 E
port 6 nsew
flabel metal3 s -24 80 -24 80 7 FreeSans 24 270 0 0 F
port 7 nsew
<< end >>
